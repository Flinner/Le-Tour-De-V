module main

fn main() {
	println('Hello!, こんにちは, مرحبا! ')
}
