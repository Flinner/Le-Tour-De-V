module main

import time

fn main() {
	println('Welcome to the playground!')

	println('The time now is $time.now()')
}
