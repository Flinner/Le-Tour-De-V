module main

fn main() {
	println('hello world!')
}

// a "hello world" program in V is as simple as

println('hello world')
