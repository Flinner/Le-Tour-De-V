// module options:

/*
*   install           Install a module from VPM.
*   remove            Remove a module that was installed from VPM.
*   search            Search for a module from VPM.
*   update            Update an installed module from VPM.
*   upgrade           Upgrade all the outdated modules.
*  list              List all installed modules.
*   outdated          Show installed modules that need updates.
*/
